CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 174 454 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
44127.9 0
0
13 Logic Switch~
5 183 370 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
44127.9 0
0
13 Logic Switch~
5 205 280 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8157 0 0
2
44127.9 0
0
13 Logic Switch~
5 207 149 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
44127.9 0
0
13 Logic Switch~
5 207 98 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
44127.9 1
0
14 Logic Display~
6 476 406 0 1 2
10 2
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
44127.9 0
0
14 Logic Display~
6 471 271 0 1 2
10 3
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
44127.9 0
0
9 Inverter~
13 344 276 0 2 22
0 7 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
972 0 0
2
44127.9 0
0
9 2-In AND~
219 346 409 0 3 22
0 6 5 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3472 0 0
2
44127.9 0
0
8 2-In OR~
219 331 118 0 3 22
0 9 8 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9998 0 0
2
5.89958e-315 0
0
14 Logic Display~
6 459 82 0 1 2
10 4
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
44127.9 2
0
8
3 1 2 0 0 8320 0 9 6 0 0 3
367 409
367 410
460 410
2 1 3 0 0 8320 0 8 7 0 0 3
365 276
365 275
455 275
1 3 4 0 0 4224 0 11 10 0 0 4
443 86
372 86
372 118
364 118
1 2 5 0 0 4224 0 1 9 0 0 4
186 454
273 454
273 418
322 418
1 1 6 0 0 4224 0 2 9 0 0 5
195 370
300 370
300 404
322 404
322 400
1 1 7 0 0 4224 0 3 8 0 0 3
217 280
329 280
329 276
1 2 8 0 0 12416 0 4 10 0 0 4
219 149
268 149
268 127
318 127
1 1 9 0 0 12416 0 5 10 0 0 4
219 98
268 98
268 109
318 109
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
